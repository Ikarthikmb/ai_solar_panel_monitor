magic
tech sky130A
magscale 1 2
timestamp 1699154466
<< obsli1 >>
rect 1104 2159 98808 597329
<< obsm1 >>
rect 934 2128 98808 597360
<< metal2 >>
rect 7194 599200 7250 600000
rect 21454 599200 21510 600000
rect 35714 599200 35770 600000
rect 49974 599200 50030 600000
rect 64234 599200 64290 600000
rect 78494 599200 78550 600000
rect 92754 599200 92810 600000
rect 10046 0 10102 800
rect 30010 0 30066 800
rect 49974 0 50030 800
rect 69938 0 69994 800
rect 89902 0 89958 800
<< obsm2 >>
rect 938 599144 7138 599298
rect 7306 599144 21398 599298
rect 21566 599144 35658 599298
rect 35826 599144 49918 599298
rect 50086 599144 64178 599298
rect 64346 599144 78438 599298
rect 78606 599144 92698 599298
rect 92866 599144 98514 599298
rect 938 856 98514 599144
rect 938 800 9990 856
rect 10158 800 29954 856
rect 30122 800 49918 856
rect 50086 800 69882 856
rect 70050 800 89846 856
rect 90014 800 98514 856
<< metal3 >>
rect 99200 584536 100000 584656
rect 0 580456 800 580576
rect 99200 559784 100000 559904
rect 0 545368 800 545488
rect 99200 535032 100000 535152
rect 0 510280 800 510400
rect 99200 510280 100000 510400
rect 99200 485528 100000 485648
rect 0 475192 800 475312
rect 99200 460776 100000 460896
rect 0 440104 800 440224
rect 99200 436024 100000 436144
rect 99200 411272 100000 411392
rect 0 405016 800 405136
rect 99200 386520 100000 386640
rect 0 369928 800 370048
rect 99200 361768 100000 361888
rect 99200 337016 100000 337136
rect 0 334840 800 334960
rect 99200 312264 100000 312384
rect 0 299752 800 299872
rect 99200 287512 100000 287632
rect 0 264664 800 264784
rect 99200 262760 100000 262880
rect 99200 238008 100000 238128
rect 0 229576 800 229696
rect 99200 213256 100000 213376
rect 0 194488 800 194608
rect 99200 188504 100000 188624
rect 99200 163752 100000 163872
rect 0 159400 800 159520
rect 99200 139000 100000 139120
rect 0 124312 800 124432
rect 99200 114248 100000 114368
rect 99200 89496 100000 89616
rect 0 89224 800 89344
rect 99200 64744 100000 64864
rect 0 54136 800 54256
rect 99200 39992 100000 40112
rect 0 19048 800 19168
rect 99200 15240 100000 15360
<< obsm3 >>
rect 798 584736 99200 597345
rect 798 584456 99120 584736
rect 798 580656 99200 584456
rect 880 580376 99200 580656
rect 798 559984 99200 580376
rect 798 559704 99120 559984
rect 798 545568 99200 559704
rect 880 545288 99200 545568
rect 798 535232 99200 545288
rect 798 534952 99120 535232
rect 798 510480 99200 534952
rect 880 510200 99120 510480
rect 798 485728 99200 510200
rect 798 485448 99120 485728
rect 798 475392 99200 485448
rect 880 475112 99200 475392
rect 798 460976 99200 475112
rect 798 460696 99120 460976
rect 798 440304 99200 460696
rect 880 440024 99200 440304
rect 798 436224 99200 440024
rect 798 435944 99120 436224
rect 798 411472 99200 435944
rect 798 411192 99120 411472
rect 798 405216 99200 411192
rect 880 404936 99200 405216
rect 798 386720 99200 404936
rect 798 386440 99120 386720
rect 798 370128 99200 386440
rect 880 369848 99200 370128
rect 798 361968 99200 369848
rect 798 361688 99120 361968
rect 798 337216 99200 361688
rect 798 336936 99120 337216
rect 798 335040 99200 336936
rect 880 334760 99200 335040
rect 798 312464 99200 334760
rect 798 312184 99120 312464
rect 798 299952 99200 312184
rect 880 299672 99200 299952
rect 798 287712 99200 299672
rect 798 287432 99120 287712
rect 798 264864 99200 287432
rect 880 264584 99200 264864
rect 798 262960 99200 264584
rect 798 262680 99120 262960
rect 798 238208 99200 262680
rect 798 237928 99120 238208
rect 798 229776 99200 237928
rect 880 229496 99200 229776
rect 798 213456 99200 229496
rect 798 213176 99120 213456
rect 798 194688 99200 213176
rect 880 194408 99200 194688
rect 798 188704 99200 194408
rect 798 188424 99120 188704
rect 798 163952 99200 188424
rect 798 163672 99120 163952
rect 798 159600 99200 163672
rect 880 159320 99200 159600
rect 798 139200 99200 159320
rect 798 138920 99120 139200
rect 798 124512 99200 138920
rect 880 124232 99200 124512
rect 798 114448 99200 124232
rect 798 114168 99120 114448
rect 798 89696 99200 114168
rect 798 89424 99120 89696
rect 880 89416 99120 89424
rect 880 89144 99200 89416
rect 798 64944 99200 89144
rect 798 64664 99120 64944
rect 798 54336 99200 64664
rect 880 54056 99200 54336
rect 798 40192 99200 54056
rect 798 39912 99120 40192
rect 798 19248 99200 39912
rect 880 18968 99200 19248
rect 798 15440 99200 18968
rect 798 15160 99120 15440
rect 798 2143 99200 15160
<< metal4 >>
rect 4208 2128 4528 597360
rect 19568 2128 19888 597360
rect 34928 2128 35248 597360
rect 50288 2128 50608 597360
rect 65648 2128 65968 597360
rect 81008 2128 81328 597360
rect 96368 2128 96688 597360
<< labels >>
rlabel metal3 s 99200 15240 100000 15360 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 369928 800 370048 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 264664 800 264784 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 0 159400 800 159520 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 0 124312 800 124432 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 0 89224 800 89344 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 0 54136 800 54256 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 92754 599200 92810 600000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 78494 599200 78550 600000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 64234 599200 64290 600000 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 99200 89496 100000 89616 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 49974 599200 50030 600000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 35714 599200 35770 600000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 21454 599200 21510 600000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 7194 599200 7250 600000 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 99200 163752 100000 163872 6 io_in[2]
port 17 nsew signal input
rlabel metal3 s 99200 238008 100000 238128 6 io_in[3]
port 18 nsew signal input
rlabel metal3 s 99200 312264 100000 312384 6 io_in[4]
port 19 nsew signal input
rlabel metal3 s 99200 386520 100000 386640 6 io_in[5]
port 20 nsew signal input
rlabel metal3 s 99200 460776 100000 460896 6 io_in[6]
port 21 nsew signal input
rlabel metal3 s 99200 535032 100000 535152 6 io_in[7]
port 22 nsew signal input
rlabel metal3 s 0 580456 800 580576 6 io_in[8]
port 23 nsew signal input
rlabel metal3 s 0 475192 800 475312 6 io_in[9]
port 24 nsew signal input
rlabel metal3 s 99200 64744 100000 64864 6 io_oeb[0]
port 25 nsew signal output
rlabel metal3 s 0 299752 800 299872 6 io_oeb[10]
port 26 nsew signal output
rlabel metal3 s 0 194488 800 194608 6 io_oeb[11]
port 27 nsew signal output
rlabel metal3 s 99200 139000 100000 139120 6 io_oeb[1]
port 28 nsew signal output
rlabel metal3 s 99200 213256 100000 213376 6 io_oeb[2]
port 29 nsew signal output
rlabel metal3 s 99200 287512 100000 287632 6 io_oeb[3]
port 30 nsew signal output
rlabel metal3 s 99200 361768 100000 361888 6 io_oeb[4]
port 31 nsew signal output
rlabel metal3 s 99200 436024 100000 436144 6 io_oeb[5]
port 32 nsew signal output
rlabel metal3 s 99200 510280 100000 510400 6 io_oeb[6]
port 33 nsew signal output
rlabel metal3 s 99200 584536 100000 584656 6 io_oeb[7]
port 34 nsew signal output
rlabel metal3 s 0 510280 800 510400 6 io_oeb[8]
port 35 nsew signal output
rlabel metal3 s 0 405016 800 405136 6 io_oeb[9]
port 36 nsew signal output
rlabel metal3 s 99200 39992 100000 40112 6 io_out[0]
port 37 nsew signal output
rlabel metal3 s 0 334840 800 334960 6 io_out[10]
port 38 nsew signal output
rlabel metal3 s 0 229576 800 229696 6 io_out[11]
port 39 nsew signal output
rlabel metal3 s 99200 114248 100000 114368 6 io_out[1]
port 40 nsew signal output
rlabel metal3 s 99200 188504 100000 188624 6 io_out[2]
port 41 nsew signal output
rlabel metal3 s 99200 262760 100000 262880 6 io_out[3]
port 42 nsew signal output
rlabel metal3 s 99200 337016 100000 337136 6 io_out[4]
port 43 nsew signal output
rlabel metal3 s 99200 411272 100000 411392 6 io_out[5]
port 44 nsew signal output
rlabel metal3 s 99200 485528 100000 485648 6 io_out[6]
port 45 nsew signal output
rlabel metal3 s 99200 559784 100000 559904 6 io_out[7]
port 46 nsew signal output
rlabel metal3 s 0 545368 800 545488 6 io_out[8]
port 47 nsew signal output
rlabel metal3 s 0 440104 800 440224 6 io_out[9]
port 48 nsew signal output
rlabel metal2 s 49974 0 50030 800 6 irq[0]
port 49 nsew signal output
rlabel metal2 s 69938 0 69994 800 6 irq[1]
port 50 nsew signal output
rlabel metal2 s 89902 0 89958 800 6 irq[2]
port 51 nsew signal output
rlabel metal4 s 4208 2128 4528 597360 6 vccd1
port 52 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 597360 6 vccd1
port 52 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 597360 6 vccd1
port 52 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 597360 6 vccd1
port 52 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 597360 6 vssd1
port 53 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 597360 6 vssd1
port 53 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 597360 6 vssd1
port 53 nsew ground bidirectional
rlabel metal2 s 10046 0 10102 800 6 wb_clk_i
port 54 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 wb_rst_i
port 55 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 100000 600000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 16128278
string GDS_FILE /Users/karthikmb/Iceberg-dir/inventory/ikarthikmb-github/ai-design-congest-oct-2023/ai_solar_panel_monitor/openlane/user_proj_solar/runs/23_11_04_22_17/results/signoff/user_proj_solar.magic.gds
string GDS_START 142108
<< end >>

