magic
tech sky130A
magscale 1 2
timestamp 1698859417
<< nwell >>
rect 1066 596485 98846 597051
rect 1066 595397 98846 595963
rect 1066 594309 98846 594875
rect 1066 593221 98846 593787
rect 1066 592133 98846 592699
rect 1066 591045 98846 591611
rect 1066 589957 98846 590523
rect 1066 588869 98846 589435
rect 1066 587781 98846 588347
rect 1066 586693 98846 587259
rect 1066 585605 98846 586171
rect 1066 584517 98846 585083
rect 1066 583429 98846 583995
rect 1066 582341 98846 582907
rect 1066 581253 98846 581819
rect 1066 580165 98846 580731
rect 1066 579077 98846 579643
rect 1066 577989 98846 578555
rect 1066 576901 98846 577467
rect 1066 575813 98846 576379
rect 1066 574725 98846 575291
rect 1066 573637 98846 574203
rect 1066 572549 98846 573115
rect 1066 571461 98846 572027
rect 1066 570373 98846 570939
rect 1066 569285 98846 569851
rect 1066 568197 98846 568763
rect 1066 567109 98846 567675
rect 1066 566021 98846 566587
rect 1066 564933 98846 565499
rect 1066 563845 98846 564411
rect 1066 562757 98846 563323
rect 1066 561669 98846 562235
rect 1066 560581 98846 561147
rect 1066 559493 98846 560059
rect 1066 558405 98846 558971
rect 1066 557317 98846 557883
rect 1066 556229 98846 556795
rect 1066 555141 98846 555707
rect 1066 554053 98846 554619
rect 1066 552965 98846 553531
rect 1066 551877 98846 552443
rect 1066 550789 98846 551355
rect 1066 549701 98846 550267
rect 1066 548613 98846 549179
rect 1066 547525 98846 548091
rect 1066 546437 98846 547003
rect 1066 545349 98846 545915
rect 1066 544261 98846 544827
rect 1066 543173 98846 543739
rect 1066 542085 98846 542651
rect 1066 540997 98846 541563
rect 1066 539909 98846 540475
rect 1066 538821 98846 539387
rect 1066 537733 98846 538299
rect 1066 536645 98846 537211
rect 1066 535557 98846 536123
rect 1066 534469 98846 535035
rect 1066 533381 98846 533947
rect 1066 532293 98846 532859
rect 1066 531205 98846 531771
rect 1066 530117 98846 530683
rect 1066 529029 98846 529595
rect 1066 527941 98846 528507
rect 1066 526853 98846 527419
rect 1066 525765 98846 526331
rect 1066 524677 98846 525243
rect 1066 523589 98846 524155
rect 1066 522501 98846 523067
rect 1066 521413 98846 521979
rect 1066 520325 98846 520891
rect 1066 519237 98846 519803
rect 1066 518149 98846 518715
rect 1066 517061 98846 517627
rect 1066 515973 98846 516539
rect 1066 514885 98846 515451
rect 1066 513797 98846 514363
rect 1066 512709 98846 513275
rect 1066 511621 98846 512187
rect 1066 510533 98846 511099
rect 1066 509445 98846 510011
rect 1066 508357 98846 508923
rect 1066 507269 98846 507835
rect 1066 506181 98846 506747
rect 1066 505093 98846 505659
rect 1066 504005 98846 504571
rect 1066 502917 98846 503483
rect 1066 501829 98846 502395
rect 1066 500741 98846 501307
rect 1066 499653 98846 500219
rect 1066 498565 98846 499131
rect 1066 497477 98846 498043
rect 1066 496389 98846 496955
rect 1066 495301 98846 495867
rect 1066 494213 98846 494779
rect 1066 493125 98846 493691
rect 1066 492037 98846 492603
rect 1066 490949 98846 491515
rect 1066 489861 98846 490427
rect 1066 488773 98846 489339
rect 1066 487685 98846 488251
rect 1066 486597 98846 487163
rect 1066 485509 98846 486075
rect 1066 484421 98846 484987
rect 1066 483333 98846 483899
rect 1066 482245 98846 482811
rect 1066 481157 98846 481723
rect 1066 480069 98846 480635
rect 1066 478981 98846 479547
rect 1066 477893 98846 478459
rect 1066 476805 98846 477371
rect 1066 475717 98846 476283
rect 1066 474629 98846 475195
rect 1066 473541 98846 474107
rect 1066 472453 98846 473019
rect 1066 471365 98846 471931
rect 1066 470277 98846 470843
rect 1066 469189 98846 469755
rect 1066 468101 98846 468667
rect 1066 467013 98846 467579
rect 1066 465925 98846 466491
rect 1066 464837 98846 465403
rect 1066 463749 98846 464315
rect 1066 462661 98846 463227
rect 1066 461573 98846 462139
rect 1066 460485 98846 461051
rect 1066 459397 98846 459963
rect 1066 458309 98846 458875
rect 1066 457221 98846 457787
rect 1066 456133 98846 456699
rect 1066 455045 98846 455611
rect 1066 453957 98846 454523
rect 1066 452869 98846 453435
rect 1066 451781 98846 452347
rect 1066 450693 98846 451259
rect 1066 449605 98846 450171
rect 1066 448517 98846 449083
rect 1066 447429 98846 447995
rect 1066 446341 98846 446907
rect 1066 445253 98846 445819
rect 1066 444165 98846 444731
rect 1066 443077 98846 443643
rect 1066 441989 98846 442555
rect 1066 440901 98846 441467
rect 1066 439813 98846 440379
rect 1066 438725 98846 439291
rect 1066 437637 98846 438203
rect 1066 436549 98846 437115
rect 1066 435461 98846 436027
rect 1066 434373 98846 434939
rect 1066 433285 98846 433851
rect 1066 432197 98846 432763
rect 1066 431109 98846 431675
rect 1066 430021 98846 430587
rect 1066 428933 98846 429499
rect 1066 427845 98846 428411
rect 1066 426757 98846 427323
rect 1066 425669 98846 426235
rect 1066 424581 98846 425147
rect 1066 423493 98846 424059
rect 1066 422405 98846 422971
rect 1066 421317 98846 421883
rect 1066 420229 98846 420795
rect 1066 419141 98846 419707
rect 1066 418053 98846 418619
rect 1066 416965 98846 417531
rect 1066 415877 98846 416443
rect 1066 414789 98846 415355
rect 1066 413701 98846 414267
rect 1066 412613 98846 413179
rect 1066 411525 98846 412091
rect 1066 410437 98846 411003
rect 1066 409349 98846 409915
rect 1066 408261 98846 408827
rect 1066 407173 98846 407739
rect 1066 406085 98846 406651
rect 1066 404997 98846 405563
rect 1066 403909 98846 404475
rect 1066 402821 98846 403387
rect 1066 401733 98846 402299
rect 1066 400645 98846 401211
rect 1066 399557 98846 400123
rect 1066 398469 98846 399035
rect 1066 397381 98846 397947
rect 1066 396293 98846 396859
rect 1066 395205 98846 395771
rect 1066 394117 98846 394683
rect 1066 393029 98846 393595
rect 1066 391941 98846 392507
rect 1066 390853 98846 391419
rect 1066 389765 98846 390331
rect 1066 388677 98846 389243
rect 1066 387589 98846 388155
rect 1066 386501 98846 387067
rect 1066 385413 98846 385979
rect 1066 384325 98846 384891
rect 1066 383237 98846 383803
rect 1066 382149 98846 382715
rect 1066 381061 98846 381627
rect 1066 379973 98846 380539
rect 1066 378885 98846 379451
rect 1066 377797 98846 378363
rect 1066 376709 98846 377275
rect 1066 375621 98846 376187
rect 1066 374533 98846 375099
rect 1066 373445 98846 374011
rect 1066 372357 98846 372923
rect 1066 371269 98846 371835
rect 1066 370181 98846 370747
rect 1066 369093 98846 369659
rect 1066 368005 98846 368571
rect 1066 366917 98846 367483
rect 1066 365829 98846 366395
rect 1066 364741 98846 365307
rect 1066 363653 98846 364219
rect 1066 362565 98846 363131
rect 1066 361477 98846 362043
rect 1066 360389 98846 360955
rect 1066 359301 98846 359867
rect 1066 358213 98846 358779
rect 1066 357125 98846 357691
rect 1066 356037 98846 356603
rect 1066 354949 98846 355515
rect 1066 353861 98846 354427
rect 1066 352773 98846 353339
rect 1066 351685 98846 352251
rect 1066 350597 98846 351163
rect 1066 349509 98846 350075
rect 1066 348421 98846 348987
rect 1066 347333 98846 347899
rect 1066 346245 98846 346811
rect 1066 345157 98846 345723
rect 1066 344069 98846 344635
rect 1066 342981 98846 343547
rect 1066 341893 98846 342459
rect 1066 340805 98846 341371
rect 1066 339717 98846 340283
rect 1066 338629 98846 339195
rect 1066 337541 98846 338107
rect 1066 336453 98846 337019
rect 1066 335365 98846 335931
rect 1066 334277 98846 334843
rect 1066 333189 98846 333755
rect 1066 332101 98846 332667
rect 1066 331013 98846 331579
rect 1066 329925 98846 330491
rect 1066 328837 98846 329403
rect 1066 327749 98846 328315
rect 1066 326661 98846 327227
rect 1066 325573 98846 326139
rect 1066 324485 98846 325051
rect 1066 323397 98846 323963
rect 1066 322309 98846 322875
rect 1066 321221 98846 321787
rect 1066 320133 98846 320699
rect 1066 319045 98846 319611
rect 1066 317957 98846 318523
rect 1066 316869 98846 317435
rect 1066 315781 98846 316347
rect 1066 314693 98846 315259
rect 1066 313605 98846 314171
rect 1066 312517 98846 313083
rect 1066 311429 98846 311995
rect 1066 310341 98846 310907
rect 1066 309253 98846 309819
rect 1066 308165 98846 308731
rect 1066 307077 98846 307643
rect 1066 305989 98846 306555
rect 1066 304901 98846 305467
rect 1066 303813 98846 304379
rect 1066 302725 98846 303291
rect 1066 301637 98846 302203
rect 1066 300549 98846 301115
rect 1066 299461 98846 300027
rect 1066 298373 98846 298939
rect 1066 297285 98846 297851
rect 1066 296197 98846 296763
rect 1066 295109 98846 295675
rect 1066 294021 98846 294587
rect 1066 292933 98846 293499
rect 1066 291845 98846 292411
rect 1066 290757 98846 291323
rect 1066 289669 98846 290235
rect 1066 288581 98846 289147
rect 1066 287493 98846 288059
rect 1066 286405 98846 286971
rect 1066 285317 98846 285883
rect 1066 284229 98846 284795
rect 1066 283141 98846 283707
rect 1066 282053 98846 282619
rect 1066 280965 98846 281531
rect 1066 279877 98846 280443
rect 1066 278789 98846 279355
rect 1066 277701 98846 278267
rect 1066 276613 98846 277179
rect 1066 275525 98846 276091
rect 1066 274437 98846 275003
rect 1066 273349 98846 273915
rect 1066 272261 98846 272827
rect 1066 271173 98846 271739
rect 1066 270085 98846 270651
rect 1066 268997 98846 269563
rect 1066 267909 98846 268475
rect 1066 266821 98846 267387
rect 1066 265733 98846 266299
rect 1066 264645 98846 265211
rect 1066 263557 98846 264123
rect 1066 262469 98846 263035
rect 1066 261381 98846 261947
rect 1066 260293 98846 260859
rect 1066 259205 98846 259771
rect 1066 258117 98846 258683
rect 1066 257029 98846 257595
rect 1066 255941 98846 256507
rect 1066 254853 98846 255419
rect 1066 253765 98846 254331
rect 1066 252677 98846 253243
rect 1066 251589 98846 252155
rect 1066 250501 98846 251067
rect 1066 249413 98846 249979
rect 1066 248325 98846 248891
rect 1066 247237 98846 247803
rect 1066 246149 98846 246715
rect 1066 245061 98846 245627
rect 1066 243973 98846 244539
rect 1066 242885 98846 243451
rect 1066 241797 98846 242363
rect 1066 240709 98846 241275
rect 1066 239621 98846 240187
rect 1066 238533 98846 239099
rect 1066 237445 98846 238011
rect 1066 236357 98846 236923
rect 1066 235269 98846 235835
rect 1066 234181 98846 234747
rect 1066 233093 98846 233659
rect 1066 232005 98846 232571
rect 1066 230917 98846 231483
rect 1066 229829 98846 230395
rect 1066 228741 98846 229307
rect 1066 227653 98846 228219
rect 1066 226565 98846 227131
rect 1066 225477 98846 226043
rect 1066 224389 98846 224955
rect 1066 223301 98846 223867
rect 1066 222213 98846 222779
rect 1066 221125 98846 221691
rect 1066 220037 98846 220603
rect 1066 218949 98846 219515
rect 1066 217861 98846 218427
rect 1066 216773 98846 217339
rect 1066 215685 98846 216251
rect 1066 214597 98846 215163
rect 1066 213509 98846 214075
rect 1066 212421 98846 212987
rect 1066 211333 98846 211899
rect 1066 210245 98846 210811
rect 1066 209157 98846 209723
rect 1066 208069 98846 208635
rect 1066 206981 98846 207547
rect 1066 205893 98846 206459
rect 1066 204805 98846 205371
rect 1066 203717 98846 204283
rect 1066 202629 98846 203195
rect 1066 201541 98846 202107
rect 1066 200453 98846 201019
rect 1066 199365 98846 199931
rect 1066 198277 98846 198843
rect 1066 197189 98846 197755
rect 1066 196101 98846 196667
rect 1066 195013 98846 195579
rect 1066 193925 98846 194491
rect 1066 192837 98846 193403
rect 1066 191749 98846 192315
rect 1066 190661 98846 191227
rect 1066 189573 98846 190139
rect 1066 188485 98846 189051
rect 1066 187397 98846 187963
rect 1066 186309 98846 186875
rect 1066 185221 98846 185787
rect 1066 184133 98846 184699
rect 1066 183045 98846 183611
rect 1066 181957 98846 182523
rect 1066 180869 98846 181435
rect 1066 179781 98846 180347
rect 1066 178693 98846 179259
rect 1066 177605 98846 178171
rect 1066 176517 98846 177083
rect 1066 175429 98846 175995
rect 1066 174341 98846 174907
rect 1066 173253 98846 173819
rect 1066 172165 98846 172731
rect 1066 171077 98846 171643
rect 1066 169989 98846 170555
rect 1066 168901 98846 169467
rect 1066 167813 98846 168379
rect 1066 166725 98846 167291
rect 1066 165637 98846 166203
rect 1066 164549 98846 165115
rect 1066 163461 98846 164027
rect 1066 162373 98846 162939
rect 1066 161285 98846 161851
rect 1066 160197 98846 160763
rect 1066 159109 98846 159675
rect 1066 158021 98846 158587
rect 1066 156933 98846 157499
rect 1066 155845 98846 156411
rect 1066 154757 98846 155323
rect 1066 153669 98846 154235
rect 1066 152581 98846 153147
rect 1066 151493 98846 152059
rect 1066 150405 98846 150971
rect 1066 149317 98846 149883
rect 1066 148229 98846 148795
rect 1066 147141 98846 147707
rect 1066 146053 98846 146619
rect 1066 144965 98846 145531
rect 1066 143877 98846 144443
rect 1066 142789 98846 143355
rect 1066 141701 98846 142267
rect 1066 140613 98846 141179
rect 1066 139525 98846 140091
rect 1066 138437 98846 139003
rect 1066 137349 98846 137915
rect 1066 136261 98846 136827
rect 1066 135173 98846 135739
rect 1066 134085 98846 134651
rect 1066 132997 98846 133563
rect 1066 131909 98846 132475
rect 1066 130821 98846 131387
rect 1066 129733 98846 130299
rect 1066 128645 98846 129211
rect 1066 127557 98846 128123
rect 1066 126469 98846 127035
rect 1066 125381 98846 125947
rect 1066 124293 98846 124859
rect 1066 123205 98846 123771
rect 1066 122117 98846 122683
rect 1066 121029 98846 121595
rect 1066 119941 98846 120507
rect 1066 118853 98846 119419
rect 1066 117765 98846 118331
rect 1066 116677 98846 117243
rect 1066 115589 98846 116155
rect 1066 114501 98846 115067
rect 1066 113413 98846 113979
rect 1066 112325 98846 112891
rect 1066 111237 98846 111803
rect 1066 110149 98846 110715
rect 1066 109061 98846 109627
rect 1066 107973 98846 108539
rect 1066 106885 98846 107451
rect 1066 105797 98846 106363
rect 1066 104709 98846 105275
rect 1066 103621 98846 104187
rect 1066 102533 98846 103099
rect 1066 101445 98846 102011
rect 1066 100357 98846 100923
rect 1066 99269 98846 99835
rect 1066 98181 98846 98747
rect 1066 97093 98846 97659
rect 1066 96005 98846 96571
rect 1066 94917 98846 95483
rect 1066 93829 98846 94395
rect 1066 92741 98846 93307
rect 1066 91653 98846 92219
rect 1066 90565 98846 91131
rect 1066 89477 98846 90043
rect 1066 88389 98846 88955
rect 1066 87301 98846 87867
rect 1066 86213 98846 86779
rect 1066 85125 98846 85691
rect 1066 84037 98846 84603
rect 1066 82949 98846 83515
rect 1066 81861 98846 82427
rect 1066 80773 98846 81339
rect 1066 79685 98846 80251
rect 1066 78597 98846 79163
rect 1066 77509 98846 78075
rect 1066 76421 98846 76987
rect 1066 75333 98846 75899
rect 1066 74245 98846 74811
rect 1066 73157 98846 73723
rect 1066 72069 98846 72635
rect 1066 70981 98846 71547
rect 1066 69893 98846 70459
rect 1066 68805 98846 69371
rect 1066 67717 98846 68283
rect 1066 66629 98846 67195
rect 1066 65541 98846 66107
rect 1066 64453 98846 65019
rect 1066 63365 98846 63931
rect 1066 62277 98846 62843
rect 1066 61189 98846 61755
rect 1066 60101 98846 60667
rect 1066 59013 98846 59579
rect 1066 57925 98846 58491
rect 1066 56837 98846 57403
rect 1066 55749 98846 56315
rect 1066 54661 98846 55227
rect 1066 53573 98846 54139
rect 1066 52485 98846 53051
rect 1066 51397 98846 51963
rect 1066 50309 98846 50875
rect 1066 49221 98846 49787
rect 1066 48133 98846 48699
rect 1066 47045 98846 47611
rect 1066 45957 98846 46523
rect 1066 44869 98846 45435
rect 1066 43781 98846 44347
rect 1066 42693 98846 43259
rect 1066 41605 98846 42171
rect 1066 40517 98846 41083
rect 1066 39429 98846 39995
rect 1066 38341 98846 38907
rect 1066 37253 98846 37819
rect 1066 36165 98846 36731
rect 1066 35077 98846 35643
rect 1066 33989 98846 34555
rect 1066 32901 98846 33467
rect 1066 31813 98846 32379
rect 1066 30725 98846 31291
rect 1066 29637 98846 30203
rect 1066 28549 98846 29115
rect 1066 27461 98846 28027
rect 1066 26373 98846 26939
rect 1066 25285 98846 25851
rect 1066 24197 98846 24763
rect 1066 23109 98846 23675
rect 1066 22021 98846 22587
rect 1066 20933 98846 21499
rect 1066 19845 98846 20411
rect 1066 18757 98846 19323
rect 1066 17669 98846 18235
rect 1066 16581 98846 17147
rect 1066 15493 98846 16059
rect 1066 14405 98846 14971
rect 1066 13317 98846 13883
rect 1066 12229 98846 12795
rect 1066 11141 98846 11707
rect 1066 10053 98846 10619
rect 1066 8965 98846 9531
rect 1066 7877 98846 8443
rect 1066 6789 98846 7355
rect 1066 5701 98846 6267
rect 1066 4613 98846 5179
rect 1066 3525 98846 4091
rect 1066 2437 98846 3003
<< obsli1 >>
rect 1104 2159 98808 597329
<< obsm1 >>
rect 1104 2128 98808 597360
<< metal2 >>
rect 2318 599200 2374 600000
rect 5722 599200 5778 600000
rect 9126 599200 9182 600000
rect 12530 599200 12586 600000
rect 15934 599200 15990 600000
rect 19338 599200 19394 600000
rect 22742 599200 22798 600000
rect 26146 599200 26202 600000
rect 29550 599200 29606 600000
rect 32954 599200 33010 600000
rect 36358 599200 36414 600000
rect 39762 599200 39818 600000
rect 43166 599200 43222 600000
rect 46570 599200 46626 600000
rect 49974 599200 50030 600000
rect 53378 599200 53434 600000
rect 56782 599200 56838 600000
rect 60186 599200 60242 600000
rect 63590 599200 63646 600000
rect 66994 599200 67050 600000
rect 70398 599200 70454 600000
rect 73802 599200 73858 600000
rect 77206 599200 77262 600000
rect 80610 599200 80666 600000
rect 84014 599200 84070 600000
rect 87418 599200 87474 600000
rect 90822 599200 90878 600000
rect 94226 599200 94282 600000
rect 97630 599200 97686 600000
rect 24950 0 25006 800
rect 74906 0 74962 800
<< obsm2 >>
rect 2430 599144 5666 599298
rect 5834 599144 9070 599298
rect 9238 599144 12474 599298
rect 12642 599144 15878 599298
rect 16046 599144 19282 599298
rect 19450 599144 22686 599298
rect 22854 599144 26090 599298
rect 26258 599144 29494 599298
rect 29662 599144 32898 599298
rect 33066 599144 36302 599298
rect 36470 599144 39706 599298
rect 39874 599144 43110 599298
rect 43278 599144 46514 599298
rect 46682 599144 49918 599298
rect 50086 599144 53322 599298
rect 53490 599144 56726 599298
rect 56894 599144 60130 599298
rect 60298 599144 63534 599298
rect 63702 599144 66938 599298
rect 67106 599144 70342 599298
rect 70510 599144 73746 599298
rect 73914 599144 77150 599298
rect 77318 599144 80554 599298
rect 80722 599144 83958 599298
rect 84126 599144 87362 599298
rect 87530 599144 90766 599298
rect 90934 599144 94170 599298
rect 94338 599144 96682 599298
rect 2374 856 96682 599144
rect 2374 800 24894 856
rect 25062 800 74850 856
rect 75018 800 96682 856
<< obsm3 >>
rect 4210 2143 96686 597345
<< metal4 >>
rect 4208 2128 4528 597360
rect 19568 2128 19888 597360
rect 34928 2128 35248 597360
rect 50288 2128 50608 597360
rect 65648 2128 65968 597360
rect 81008 2128 81328 597360
rect 96368 2128 96688 597360
<< labels >>
rlabel metal2 s 97630 599200 97686 600000 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 63590 599200 63646 600000 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 60186 599200 60242 600000 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 56782 599200 56838 600000 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 53378 599200 53434 600000 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 49974 599200 50030 600000 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 46570 599200 46626 600000 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 43166 599200 43222 600000 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal2 s 39762 599200 39818 600000 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal2 s 36358 599200 36414 600000 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal2 s 32954 599200 33010 600000 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal2 s 94226 599200 94282 600000 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal2 s 29550 599200 29606 600000 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal2 s 26146 599200 26202 600000 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal2 s 22742 599200 22798 600000 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal2 s 19338 599200 19394 600000 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal2 s 15934 599200 15990 600000 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal2 s 12530 599200 12586 600000 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal2 s 9126 599200 9182 600000 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal2 s 5722 599200 5778 600000 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal2 s 2318 599200 2374 600000 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal2 s 90822 599200 90878 600000 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal2 s 87418 599200 87474 600000 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal2 s 84014 599200 84070 600000 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal2 s 80610 599200 80666 600000 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal2 s 77206 599200 77262 600000 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal2 s 73802 599200 73858 600000 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 70398 599200 70454 600000 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 66994 599200 67050 600000 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal4 s 4208 2128 4528 597360 6 vccd1
port 30 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 597360 6 vccd1
port 30 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 597360 6 vccd1
port 30 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 597360 6 vccd1
port 30 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 597360 6 vssd1
port 31 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 597360 6 vssd1
port 31 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 597360 6 vssd1
port 31 nsew ground bidirectional
rlabel metal2 s 24950 0 25006 800 6 wb_clk_i
port 32 nsew signal input
rlabel metal2 s 74906 0 74962 800 6 wb_rst_i
port 33 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 100000 600000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 15844046
string GDS_FILE /Users/karthikmb/Iceberg-dir/inventory/ikarthikmb-github/ai-design-congest-oct-2023/ai_solar_panel_monitor/openlane/user_proj_solar/runs/23_11_01_12_20/results/signoff/user_proj_solar.magic.gds
string GDS_START 94086
<< end >>

