VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_solar
  CLASS BLOCK ;
  FOREIGN user_proj_solar ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 3000.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 76.200 500.000 76.800 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1849.640 4.000 1850.240 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1323.320 4.000 1323.920 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 797.000 4.000 797.600 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 621.560 4.000 622.160 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.120 4.000 446.720 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 2996.000 464.050 3000.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.470 2996.000 392.750 3000.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 2996.000 321.450 3000.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 447.480 500.000 448.080 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 2996.000 250.150 3000.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 2996.000 178.850 3000.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 2996.000 107.550 3000.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 2996.000 36.250 3000.000 ;
    END
  END io_in[23]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 818.760 500.000 819.360 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 1190.040 500.000 1190.640 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 1561.320 500.000 1561.920 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 1932.600 500.000 1933.200 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 2303.880 500.000 2304.480 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 2675.160 500.000 2675.760 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2902.280 4.000 2902.880 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2375.960 4.000 2376.560 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 323.720 500.000 324.320 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1498.760 4.000 1499.360 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 972.440 4.000 973.040 ;
    END
  END io_oeb[11]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 695.000 500.000 695.600 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 1066.280 500.000 1066.880 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 1437.560 500.000 1438.160 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 1808.840 500.000 1809.440 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 2180.120 500.000 2180.720 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 2551.400 500.000 2552.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 2922.680 500.000 2923.280 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2551.400 4.000 2552.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2025.080 4.000 2025.680 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 199.960 500.000 200.560 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1674.200 4.000 1674.800 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1147.880 4.000 1148.480 ;
    END
  END io_out[11]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 571.240 500.000 571.840 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 942.520 500.000 943.120 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 1313.800 500.000 1314.400 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 1685.080 500.000 1685.680 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 2056.360 500.000 2056.960 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 2427.640 500.000 2428.240 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 2798.920 500.000 2799.520 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2726.840 4.000 2727.440 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2200.520 4.000 2201.120 ;
    END
  END io_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 2986.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 2986.800 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END wb_rst_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 494.040 2986.645 ;
      LAYER met1 ;
        RECT 4.670 10.640 494.430 2986.800 ;
      LAYER met2 ;
        RECT 4.690 4.280 494.410 2986.745 ;
        RECT 4.690 4.000 124.470 4.280 ;
        RECT 125.310 4.000 374.250 4.280 ;
        RECT 375.090 4.000 494.410 4.280 ;
      LAYER met3 ;
        RECT 3.990 2923.680 496.000 2986.725 ;
        RECT 3.990 2922.280 495.600 2923.680 ;
        RECT 3.990 2903.280 496.000 2922.280 ;
        RECT 4.400 2901.880 496.000 2903.280 ;
        RECT 3.990 2799.920 496.000 2901.880 ;
        RECT 3.990 2798.520 495.600 2799.920 ;
        RECT 3.990 2727.840 496.000 2798.520 ;
        RECT 4.400 2726.440 496.000 2727.840 ;
        RECT 3.990 2676.160 496.000 2726.440 ;
        RECT 3.990 2674.760 495.600 2676.160 ;
        RECT 3.990 2552.400 496.000 2674.760 ;
        RECT 4.400 2551.000 495.600 2552.400 ;
        RECT 3.990 2428.640 496.000 2551.000 ;
        RECT 3.990 2427.240 495.600 2428.640 ;
        RECT 3.990 2376.960 496.000 2427.240 ;
        RECT 4.400 2375.560 496.000 2376.960 ;
        RECT 3.990 2304.880 496.000 2375.560 ;
        RECT 3.990 2303.480 495.600 2304.880 ;
        RECT 3.990 2201.520 496.000 2303.480 ;
        RECT 4.400 2200.120 496.000 2201.520 ;
        RECT 3.990 2181.120 496.000 2200.120 ;
        RECT 3.990 2179.720 495.600 2181.120 ;
        RECT 3.990 2057.360 496.000 2179.720 ;
        RECT 3.990 2055.960 495.600 2057.360 ;
        RECT 3.990 2026.080 496.000 2055.960 ;
        RECT 4.400 2024.680 496.000 2026.080 ;
        RECT 3.990 1933.600 496.000 2024.680 ;
        RECT 3.990 1932.200 495.600 1933.600 ;
        RECT 3.990 1850.640 496.000 1932.200 ;
        RECT 4.400 1849.240 496.000 1850.640 ;
        RECT 3.990 1809.840 496.000 1849.240 ;
        RECT 3.990 1808.440 495.600 1809.840 ;
        RECT 3.990 1686.080 496.000 1808.440 ;
        RECT 3.990 1684.680 495.600 1686.080 ;
        RECT 3.990 1675.200 496.000 1684.680 ;
        RECT 4.400 1673.800 496.000 1675.200 ;
        RECT 3.990 1562.320 496.000 1673.800 ;
        RECT 3.990 1560.920 495.600 1562.320 ;
        RECT 3.990 1499.760 496.000 1560.920 ;
        RECT 4.400 1498.360 496.000 1499.760 ;
        RECT 3.990 1438.560 496.000 1498.360 ;
        RECT 3.990 1437.160 495.600 1438.560 ;
        RECT 3.990 1324.320 496.000 1437.160 ;
        RECT 4.400 1322.920 496.000 1324.320 ;
        RECT 3.990 1314.800 496.000 1322.920 ;
        RECT 3.990 1313.400 495.600 1314.800 ;
        RECT 3.990 1191.040 496.000 1313.400 ;
        RECT 3.990 1189.640 495.600 1191.040 ;
        RECT 3.990 1148.880 496.000 1189.640 ;
        RECT 4.400 1147.480 496.000 1148.880 ;
        RECT 3.990 1067.280 496.000 1147.480 ;
        RECT 3.990 1065.880 495.600 1067.280 ;
        RECT 3.990 973.440 496.000 1065.880 ;
        RECT 4.400 972.040 496.000 973.440 ;
        RECT 3.990 943.520 496.000 972.040 ;
        RECT 3.990 942.120 495.600 943.520 ;
        RECT 3.990 819.760 496.000 942.120 ;
        RECT 3.990 818.360 495.600 819.760 ;
        RECT 3.990 798.000 496.000 818.360 ;
        RECT 4.400 796.600 496.000 798.000 ;
        RECT 3.990 696.000 496.000 796.600 ;
        RECT 3.990 694.600 495.600 696.000 ;
        RECT 3.990 622.560 496.000 694.600 ;
        RECT 4.400 621.160 496.000 622.560 ;
        RECT 3.990 572.240 496.000 621.160 ;
        RECT 3.990 570.840 495.600 572.240 ;
        RECT 3.990 448.480 496.000 570.840 ;
        RECT 3.990 447.120 495.600 448.480 ;
        RECT 4.400 447.080 495.600 447.120 ;
        RECT 4.400 445.720 496.000 447.080 ;
        RECT 3.990 324.720 496.000 445.720 ;
        RECT 3.990 323.320 495.600 324.720 ;
        RECT 3.990 271.680 496.000 323.320 ;
        RECT 4.400 270.280 496.000 271.680 ;
        RECT 3.990 200.960 496.000 270.280 ;
        RECT 3.990 199.560 495.600 200.960 ;
        RECT 3.990 96.240 496.000 199.560 ;
        RECT 4.400 94.840 496.000 96.240 ;
        RECT 3.990 77.200 496.000 94.840 ;
        RECT 3.990 75.800 495.600 77.200 ;
        RECT 3.990 10.715 496.000 75.800 ;
  END
END user_proj_solar
END LIBRARY

