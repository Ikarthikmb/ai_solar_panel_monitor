VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_solar
  CLASS BLOCK ;
  FOREIGN user_proj_solar ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 3000.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.150 2996.000 488.430 3000.000 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 2996.000 318.230 3000.000 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 2996.000 301.210 3000.000 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 283.910 2996.000 284.190 3000.000 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 266.890 2996.000 267.170 3000.000 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 249.870 2996.000 250.150 3000.000 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 232.850 2996.000 233.130 3000.000 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 215.830 2996.000 216.110 3000.000 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 198.810 2996.000 199.090 3000.000 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 181.790 2996.000 182.070 3000.000 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 164.770 2996.000 165.050 3000.000 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.130 2996.000 471.410 3000.000 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 147.750 2996.000 148.030 3000.000 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 130.730 2996.000 131.010 3000.000 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 2996.000 113.990 3000.000 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 2996.000 96.970 3000.000 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 2996.000 79.950 3000.000 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 2996.000 62.930 3000.000 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 2996.000 45.910 3000.000 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 2996.000 28.890 3000.000 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 2996.000 11.870 3000.000 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 2996.000 454.390 3000.000 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 2996.000 437.370 3000.000 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.070 2996.000 420.350 3000.000 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.050 2996.000 403.330 3000.000 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 2996.000 386.310 3000.000 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.010 2996.000 369.290 3000.000 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 2996.000 352.270 3000.000 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 2996.000 335.250 3000.000 ;
    END
  END analog_io[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 2986.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 2986.800 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END wb_rst_i
  OBS
      LAYER nwell ;
        RECT 5.330 2982.425 494.230 2985.255 ;
        RECT 5.330 2976.985 494.230 2979.815 ;
        RECT 5.330 2971.545 494.230 2974.375 ;
        RECT 5.330 2966.105 494.230 2968.935 ;
        RECT 5.330 2960.665 494.230 2963.495 ;
        RECT 5.330 2955.225 494.230 2958.055 ;
        RECT 5.330 2949.785 494.230 2952.615 ;
        RECT 5.330 2944.345 494.230 2947.175 ;
        RECT 5.330 2938.905 494.230 2941.735 ;
        RECT 5.330 2933.465 494.230 2936.295 ;
        RECT 5.330 2928.025 494.230 2930.855 ;
        RECT 5.330 2922.585 494.230 2925.415 ;
        RECT 5.330 2917.145 494.230 2919.975 ;
        RECT 5.330 2911.705 494.230 2914.535 ;
        RECT 5.330 2906.265 494.230 2909.095 ;
        RECT 5.330 2900.825 494.230 2903.655 ;
        RECT 5.330 2895.385 494.230 2898.215 ;
        RECT 5.330 2889.945 494.230 2892.775 ;
        RECT 5.330 2884.505 494.230 2887.335 ;
        RECT 5.330 2879.065 494.230 2881.895 ;
        RECT 5.330 2873.625 494.230 2876.455 ;
        RECT 5.330 2868.185 494.230 2871.015 ;
        RECT 5.330 2862.745 494.230 2865.575 ;
        RECT 5.330 2857.305 494.230 2860.135 ;
        RECT 5.330 2851.865 494.230 2854.695 ;
        RECT 5.330 2846.425 494.230 2849.255 ;
        RECT 5.330 2840.985 494.230 2843.815 ;
        RECT 5.330 2835.545 494.230 2838.375 ;
        RECT 5.330 2830.105 494.230 2832.935 ;
        RECT 5.330 2824.665 494.230 2827.495 ;
        RECT 5.330 2819.225 494.230 2822.055 ;
        RECT 5.330 2813.785 494.230 2816.615 ;
        RECT 5.330 2808.345 494.230 2811.175 ;
        RECT 5.330 2802.905 494.230 2805.735 ;
        RECT 5.330 2797.465 494.230 2800.295 ;
        RECT 5.330 2792.025 494.230 2794.855 ;
        RECT 5.330 2786.585 494.230 2789.415 ;
        RECT 5.330 2781.145 494.230 2783.975 ;
        RECT 5.330 2775.705 494.230 2778.535 ;
        RECT 5.330 2770.265 494.230 2773.095 ;
        RECT 5.330 2764.825 494.230 2767.655 ;
        RECT 5.330 2759.385 494.230 2762.215 ;
        RECT 5.330 2753.945 494.230 2756.775 ;
        RECT 5.330 2748.505 494.230 2751.335 ;
        RECT 5.330 2743.065 494.230 2745.895 ;
        RECT 5.330 2737.625 494.230 2740.455 ;
        RECT 5.330 2732.185 494.230 2735.015 ;
        RECT 5.330 2726.745 494.230 2729.575 ;
        RECT 5.330 2721.305 494.230 2724.135 ;
        RECT 5.330 2715.865 494.230 2718.695 ;
        RECT 5.330 2710.425 494.230 2713.255 ;
        RECT 5.330 2704.985 494.230 2707.815 ;
        RECT 5.330 2699.545 494.230 2702.375 ;
        RECT 5.330 2694.105 494.230 2696.935 ;
        RECT 5.330 2688.665 494.230 2691.495 ;
        RECT 5.330 2683.225 494.230 2686.055 ;
        RECT 5.330 2677.785 494.230 2680.615 ;
        RECT 5.330 2672.345 494.230 2675.175 ;
        RECT 5.330 2666.905 494.230 2669.735 ;
        RECT 5.330 2661.465 494.230 2664.295 ;
        RECT 5.330 2656.025 494.230 2658.855 ;
        RECT 5.330 2650.585 494.230 2653.415 ;
        RECT 5.330 2645.145 494.230 2647.975 ;
        RECT 5.330 2639.705 494.230 2642.535 ;
        RECT 5.330 2634.265 494.230 2637.095 ;
        RECT 5.330 2628.825 494.230 2631.655 ;
        RECT 5.330 2623.385 494.230 2626.215 ;
        RECT 5.330 2617.945 494.230 2620.775 ;
        RECT 5.330 2612.505 494.230 2615.335 ;
        RECT 5.330 2607.065 494.230 2609.895 ;
        RECT 5.330 2601.625 494.230 2604.455 ;
        RECT 5.330 2596.185 494.230 2599.015 ;
        RECT 5.330 2590.745 494.230 2593.575 ;
        RECT 5.330 2585.305 494.230 2588.135 ;
        RECT 5.330 2579.865 494.230 2582.695 ;
        RECT 5.330 2574.425 494.230 2577.255 ;
        RECT 5.330 2568.985 494.230 2571.815 ;
        RECT 5.330 2563.545 494.230 2566.375 ;
        RECT 5.330 2558.105 494.230 2560.935 ;
        RECT 5.330 2552.665 494.230 2555.495 ;
        RECT 5.330 2547.225 494.230 2550.055 ;
        RECT 5.330 2541.785 494.230 2544.615 ;
        RECT 5.330 2536.345 494.230 2539.175 ;
        RECT 5.330 2530.905 494.230 2533.735 ;
        RECT 5.330 2525.465 494.230 2528.295 ;
        RECT 5.330 2520.025 494.230 2522.855 ;
        RECT 5.330 2514.585 494.230 2517.415 ;
        RECT 5.330 2509.145 494.230 2511.975 ;
        RECT 5.330 2503.705 494.230 2506.535 ;
        RECT 5.330 2498.265 494.230 2501.095 ;
        RECT 5.330 2492.825 494.230 2495.655 ;
        RECT 5.330 2487.385 494.230 2490.215 ;
        RECT 5.330 2481.945 494.230 2484.775 ;
        RECT 5.330 2476.505 494.230 2479.335 ;
        RECT 5.330 2471.065 494.230 2473.895 ;
        RECT 5.330 2465.625 494.230 2468.455 ;
        RECT 5.330 2460.185 494.230 2463.015 ;
        RECT 5.330 2454.745 494.230 2457.575 ;
        RECT 5.330 2449.305 494.230 2452.135 ;
        RECT 5.330 2443.865 494.230 2446.695 ;
        RECT 5.330 2438.425 494.230 2441.255 ;
        RECT 5.330 2432.985 494.230 2435.815 ;
        RECT 5.330 2427.545 494.230 2430.375 ;
        RECT 5.330 2422.105 494.230 2424.935 ;
        RECT 5.330 2416.665 494.230 2419.495 ;
        RECT 5.330 2411.225 494.230 2414.055 ;
        RECT 5.330 2405.785 494.230 2408.615 ;
        RECT 5.330 2400.345 494.230 2403.175 ;
        RECT 5.330 2394.905 494.230 2397.735 ;
        RECT 5.330 2389.465 494.230 2392.295 ;
        RECT 5.330 2384.025 494.230 2386.855 ;
        RECT 5.330 2378.585 494.230 2381.415 ;
        RECT 5.330 2373.145 494.230 2375.975 ;
        RECT 5.330 2367.705 494.230 2370.535 ;
        RECT 5.330 2362.265 494.230 2365.095 ;
        RECT 5.330 2356.825 494.230 2359.655 ;
        RECT 5.330 2351.385 494.230 2354.215 ;
        RECT 5.330 2345.945 494.230 2348.775 ;
        RECT 5.330 2340.505 494.230 2343.335 ;
        RECT 5.330 2335.065 494.230 2337.895 ;
        RECT 5.330 2329.625 494.230 2332.455 ;
        RECT 5.330 2324.185 494.230 2327.015 ;
        RECT 5.330 2318.745 494.230 2321.575 ;
        RECT 5.330 2313.305 494.230 2316.135 ;
        RECT 5.330 2307.865 494.230 2310.695 ;
        RECT 5.330 2302.425 494.230 2305.255 ;
        RECT 5.330 2296.985 494.230 2299.815 ;
        RECT 5.330 2291.545 494.230 2294.375 ;
        RECT 5.330 2286.105 494.230 2288.935 ;
        RECT 5.330 2280.665 494.230 2283.495 ;
        RECT 5.330 2275.225 494.230 2278.055 ;
        RECT 5.330 2269.785 494.230 2272.615 ;
        RECT 5.330 2264.345 494.230 2267.175 ;
        RECT 5.330 2258.905 494.230 2261.735 ;
        RECT 5.330 2253.465 494.230 2256.295 ;
        RECT 5.330 2248.025 494.230 2250.855 ;
        RECT 5.330 2242.585 494.230 2245.415 ;
        RECT 5.330 2237.145 494.230 2239.975 ;
        RECT 5.330 2231.705 494.230 2234.535 ;
        RECT 5.330 2226.265 494.230 2229.095 ;
        RECT 5.330 2220.825 494.230 2223.655 ;
        RECT 5.330 2215.385 494.230 2218.215 ;
        RECT 5.330 2209.945 494.230 2212.775 ;
        RECT 5.330 2204.505 494.230 2207.335 ;
        RECT 5.330 2199.065 494.230 2201.895 ;
        RECT 5.330 2193.625 494.230 2196.455 ;
        RECT 5.330 2188.185 494.230 2191.015 ;
        RECT 5.330 2182.745 494.230 2185.575 ;
        RECT 5.330 2177.305 494.230 2180.135 ;
        RECT 5.330 2171.865 494.230 2174.695 ;
        RECT 5.330 2166.425 494.230 2169.255 ;
        RECT 5.330 2160.985 494.230 2163.815 ;
        RECT 5.330 2155.545 494.230 2158.375 ;
        RECT 5.330 2150.105 494.230 2152.935 ;
        RECT 5.330 2144.665 494.230 2147.495 ;
        RECT 5.330 2139.225 494.230 2142.055 ;
        RECT 5.330 2133.785 494.230 2136.615 ;
        RECT 5.330 2128.345 494.230 2131.175 ;
        RECT 5.330 2122.905 494.230 2125.735 ;
        RECT 5.330 2117.465 494.230 2120.295 ;
        RECT 5.330 2112.025 494.230 2114.855 ;
        RECT 5.330 2106.585 494.230 2109.415 ;
        RECT 5.330 2101.145 494.230 2103.975 ;
        RECT 5.330 2095.705 494.230 2098.535 ;
        RECT 5.330 2090.265 494.230 2093.095 ;
        RECT 5.330 2084.825 494.230 2087.655 ;
        RECT 5.330 2079.385 494.230 2082.215 ;
        RECT 5.330 2073.945 494.230 2076.775 ;
        RECT 5.330 2068.505 494.230 2071.335 ;
        RECT 5.330 2063.065 494.230 2065.895 ;
        RECT 5.330 2057.625 494.230 2060.455 ;
        RECT 5.330 2052.185 494.230 2055.015 ;
        RECT 5.330 2046.745 494.230 2049.575 ;
        RECT 5.330 2041.305 494.230 2044.135 ;
        RECT 5.330 2035.865 494.230 2038.695 ;
        RECT 5.330 2030.425 494.230 2033.255 ;
        RECT 5.330 2024.985 494.230 2027.815 ;
        RECT 5.330 2019.545 494.230 2022.375 ;
        RECT 5.330 2014.105 494.230 2016.935 ;
        RECT 5.330 2008.665 494.230 2011.495 ;
        RECT 5.330 2003.225 494.230 2006.055 ;
        RECT 5.330 1997.785 494.230 2000.615 ;
        RECT 5.330 1992.345 494.230 1995.175 ;
        RECT 5.330 1986.905 494.230 1989.735 ;
        RECT 5.330 1981.465 494.230 1984.295 ;
        RECT 5.330 1976.025 494.230 1978.855 ;
        RECT 5.330 1970.585 494.230 1973.415 ;
        RECT 5.330 1965.145 494.230 1967.975 ;
        RECT 5.330 1959.705 494.230 1962.535 ;
        RECT 5.330 1954.265 494.230 1957.095 ;
        RECT 5.330 1948.825 494.230 1951.655 ;
        RECT 5.330 1943.385 494.230 1946.215 ;
        RECT 5.330 1937.945 494.230 1940.775 ;
        RECT 5.330 1932.505 494.230 1935.335 ;
        RECT 5.330 1927.065 494.230 1929.895 ;
        RECT 5.330 1921.625 494.230 1924.455 ;
        RECT 5.330 1916.185 494.230 1919.015 ;
        RECT 5.330 1910.745 494.230 1913.575 ;
        RECT 5.330 1905.305 494.230 1908.135 ;
        RECT 5.330 1899.865 494.230 1902.695 ;
        RECT 5.330 1894.425 494.230 1897.255 ;
        RECT 5.330 1888.985 494.230 1891.815 ;
        RECT 5.330 1883.545 494.230 1886.375 ;
        RECT 5.330 1878.105 494.230 1880.935 ;
        RECT 5.330 1872.665 494.230 1875.495 ;
        RECT 5.330 1867.225 494.230 1870.055 ;
        RECT 5.330 1861.785 494.230 1864.615 ;
        RECT 5.330 1856.345 494.230 1859.175 ;
        RECT 5.330 1850.905 494.230 1853.735 ;
        RECT 5.330 1845.465 494.230 1848.295 ;
        RECT 5.330 1840.025 494.230 1842.855 ;
        RECT 5.330 1834.585 494.230 1837.415 ;
        RECT 5.330 1829.145 494.230 1831.975 ;
        RECT 5.330 1823.705 494.230 1826.535 ;
        RECT 5.330 1818.265 494.230 1821.095 ;
        RECT 5.330 1812.825 494.230 1815.655 ;
        RECT 5.330 1807.385 494.230 1810.215 ;
        RECT 5.330 1801.945 494.230 1804.775 ;
        RECT 5.330 1796.505 494.230 1799.335 ;
        RECT 5.330 1791.065 494.230 1793.895 ;
        RECT 5.330 1785.625 494.230 1788.455 ;
        RECT 5.330 1780.185 494.230 1783.015 ;
        RECT 5.330 1774.745 494.230 1777.575 ;
        RECT 5.330 1769.305 494.230 1772.135 ;
        RECT 5.330 1763.865 494.230 1766.695 ;
        RECT 5.330 1758.425 494.230 1761.255 ;
        RECT 5.330 1752.985 494.230 1755.815 ;
        RECT 5.330 1747.545 494.230 1750.375 ;
        RECT 5.330 1742.105 494.230 1744.935 ;
        RECT 5.330 1736.665 494.230 1739.495 ;
        RECT 5.330 1731.225 494.230 1734.055 ;
        RECT 5.330 1725.785 494.230 1728.615 ;
        RECT 5.330 1720.345 494.230 1723.175 ;
        RECT 5.330 1714.905 494.230 1717.735 ;
        RECT 5.330 1709.465 494.230 1712.295 ;
        RECT 5.330 1704.025 494.230 1706.855 ;
        RECT 5.330 1698.585 494.230 1701.415 ;
        RECT 5.330 1693.145 494.230 1695.975 ;
        RECT 5.330 1687.705 494.230 1690.535 ;
        RECT 5.330 1682.265 494.230 1685.095 ;
        RECT 5.330 1676.825 494.230 1679.655 ;
        RECT 5.330 1671.385 494.230 1674.215 ;
        RECT 5.330 1665.945 494.230 1668.775 ;
        RECT 5.330 1660.505 494.230 1663.335 ;
        RECT 5.330 1655.065 494.230 1657.895 ;
        RECT 5.330 1649.625 494.230 1652.455 ;
        RECT 5.330 1644.185 494.230 1647.015 ;
        RECT 5.330 1638.745 494.230 1641.575 ;
        RECT 5.330 1633.305 494.230 1636.135 ;
        RECT 5.330 1627.865 494.230 1630.695 ;
        RECT 5.330 1622.425 494.230 1625.255 ;
        RECT 5.330 1616.985 494.230 1619.815 ;
        RECT 5.330 1611.545 494.230 1614.375 ;
        RECT 5.330 1606.105 494.230 1608.935 ;
        RECT 5.330 1600.665 494.230 1603.495 ;
        RECT 5.330 1595.225 494.230 1598.055 ;
        RECT 5.330 1589.785 494.230 1592.615 ;
        RECT 5.330 1584.345 494.230 1587.175 ;
        RECT 5.330 1578.905 494.230 1581.735 ;
        RECT 5.330 1573.465 494.230 1576.295 ;
        RECT 5.330 1568.025 494.230 1570.855 ;
        RECT 5.330 1562.585 494.230 1565.415 ;
        RECT 5.330 1557.145 494.230 1559.975 ;
        RECT 5.330 1551.705 494.230 1554.535 ;
        RECT 5.330 1546.265 494.230 1549.095 ;
        RECT 5.330 1540.825 494.230 1543.655 ;
        RECT 5.330 1535.385 494.230 1538.215 ;
        RECT 5.330 1529.945 494.230 1532.775 ;
        RECT 5.330 1524.505 494.230 1527.335 ;
        RECT 5.330 1519.065 494.230 1521.895 ;
        RECT 5.330 1513.625 494.230 1516.455 ;
        RECT 5.330 1508.185 494.230 1511.015 ;
        RECT 5.330 1502.745 494.230 1505.575 ;
        RECT 5.330 1497.305 494.230 1500.135 ;
        RECT 5.330 1491.865 494.230 1494.695 ;
        RECT 5.330 1486.425 494.230 1489.255 ;
        RECT 5.330 1480.985 494.230 1483.815 ;
        RECT 5.330 1475.545 494.230 1478.375 ;
        RECT 5.330 1470.105 494.230 1472.935 ;
        RECT 5.330 1464.665 494.230 1467.495 ;
        RECT 5.330 1459.225 494.230 1462.055 ;
        RECT 5.330 1453.785 494.230 1456.615 ;
        RECT 5.330 1448.345 494.230 1451.175 ;
        RECT 5.330 1442.905 494.230 1445.735 ;
        RECT 5.330 1437.465 494.230 1440.295 ;
        RECT 5.330 1432.025 494.230 1434.855 ;
        RECT 5.330 1426.585 494.230 1429.415 ;
        RECT 5.330 1421.145 494.230 1423.975 ;
        RECT 5.330 1415.705 494.230 1418.535 ;
        RECT 5.330 1410.265 494.230 1413.095 ;
        RECT 5.330 1404.825 494.230 1407.655 ;
        RECT 5.330 1399.385 494.230 1402.215 ;
        RECT 5.330 1393.945 494.230 1396.775 ;
        RECT 5.330 1388.505 494.230 1391.335 ;
        RECT 5.330 1383.065 494.230 1385.895 ;
        RECT 5.330 1377.625 494.230 1380.455 ;
        RECT 5.330 1372.185 494.230 1375.015 ;
        RECT 5.330 1366.745 494.230 1369.575 ;
        RECT 5.330 1361.305 494.230 1364.135 ;
        RECT 5.330 1355.865 494.230 1358.695 ;
        RECT 5.330 1350.425 494.230 1353.255 ;
        RECT 5.330 1344.985 494.230 1347.815 ;
        RECT 5.330 1339.545 494.230 1342.375 ;
        RECT 5.330 1334.105 494.230 1336.935 ;
        RECT 5.330 1328.665 494.230 1331.495 ;
        RECT 5.330 1323.225 494.230 1326.055 ;
        RECT 5.330 1317.785 494.230 1320.615 ;
        RECT 5.330 1312.345 494.230 1315.175 ;
        RECT 5.330 1306.905 494.230 1309.735 ;
        RECT 5.330 1301.465 494.230 1304.295 ;
        RECT 5.330 1296.025 494.230 1298.855 ;
        RECT 5.330 1290.585 494.230 1293.415 ;
        RECT 5.330 1285.145 494.230 1287.975 ;
        RECT 5.330 1279.705 494.230 1282.535 ;
        RECT 5.330 1274.265 494.230 1277.095 ;
        RECT 5.330 1268.825 494.230 1271.655 ;
        RECT 5.330 1263.385 494.230 1266.215 ;
        RECT 5.330 1257.945 494.230 1260.775 ;
        RECT 5.330 1252.505 494.230 1255.335 ;
        RECT 5.330 1247.065 494.230 1249.895 ;
        RECT 5.330 1241.625 494.230 1244.455 ;
        RECT 5.330 1236.185 494.230 1239.015 ;
        RECT 5.330 1230.745 494.230 1233.575 ;
        RECT 5.330 1225.305 494.230 1228.135 ;
        RECT 5.330 1219.865 494.230 1222.695 ;
        RECT 5.330 1214.425 494.230 1217.255 ;
        RECT 5.330 1208.985 494.230 1211.815 ;
        RECT 5.330 1203.545 494.230 1206.375 ;
        RECT 5.330 1198.105 494.230 1200.935 ;
        RECT 5.330 1192.665 494.230 1195.495 ;
        RECT 5.330 1187.225 494.230 1190.055 ;
        RECT 5.330 1181.785 494.230 1184.615 ;
        RECT 5.330 1176.345 494.230 1179.175 ;
        RECT 5.330 1170.905 494.230 1173.735 ;
        RECT 5.330 1165.465 494.230 1168.295 ;
        RECT 5.330 1160.025 494.230 1162.855 ;
        RECT 5.330 1154.585 494.230 1157.415 ;
        RECT 5.330 1149.145 494.230 1151.975 ;
        RECT 5.330 1143.705 494.230 1146.535 ;
        RECT 5.330 1138.265 494.230 1141.095 ;
        RECT 5.330 1132.825 494.230 1135.655 ;
        RECT 5.330 1127.385 494.230 1130.215 ;
        RECT 5.330 1121.945 494.230 1124.775 ;
        RECT 5.330 1116.505 494.230 1119.335 ;
        RECT 5.330 1111.065 494.230 1113.895 ;
        RECT 5.330 1105.625 494.230 1108.455 ;
        RECT 5.330 1100.185 494.230 1103.015 ;
        RECT 5.330 1094.745 494.230 1097.575 ;
        RECT 5.330 1089.305 494.230 1092.135 ;
        RECT 5.330 1083.865 494.230 1086.695 ;
        RECT 5.330 1078.425 494.230 1081.255 ;
        RECT 5.330 1072.985 494.230 1075.815 ;
        RECT 5.330 1067.545 494.230 1070.375 ;
        RECT 5.330 1062.105 494.230 1064.935 ;
        RECT 5.330 1056.665 494.230 1059.495 ;
        RECT 5.330 1051.225 494.230 1054.055 ;
        RECT 5.330 1045.785 494.230 1048.615 ;
        RECT 5.330 1040.345 494.230 1043.175 ;
        RECT 5.330 1034.905 494.230 1037.735 ;
        RECT 5.330 1029.465 494.230 1032.295 ;
        RECT 5.330 1024.025 494.230 1026.855 ;
        RECT 5.330 1018.585 494.230 1021.415 ;
        RECT 5.330 1013.145 494.230 1015.975 ;
        RECT 5.330 1007.705 494.230 1010.535 ;
        RECT 5.330 1002.265 494.230 1005.095 ;
        RECT 5.330 996.825 494.230 999.655 ;
        RECT 5.330 991.385 494.230 994.215 ;
        RECT 5.330 985.945 494.230 988.775 ;
        RECT 5.330 980.505 494.230 983.335 ;
        RECT 5.330 975.065 494.230 977.895 ;
        RECT 5.330 969.625 494.230 972.455 ;
        RECT 5.330 964.185 494.230 967.015 ;
        RECT 5.330 958.745 494.230 961.575 ;
        RECT 5.330 953.305 494.230 956.135 ;
        RECT 5.330 947.865 494.230 950.695 ;
        RECT 5.330 942.425 494.230 945.255 ;
        RECT 5.330 936.985 494.230 939.815 ;
        RECT 5.330 931.545 494.230 934.375 ;
        RECT 5.330 926.105 494.230 928.935 ;
        RECT 5.330 920.665 494.230 923.495 ;
        RECT 5.330 915.225 494.230 918.055 ;
        RECT 5.330 909.785 494.230 912.615 ;
        RECT 5.330 904.345 494.230 907.175 ;
        RECT 5.330 898.905 494.230 901.735 ;
        RECT 5.330 893.465 494.230 896.295 ;
        RECT 5.330 888.025 494.230 890.855 ;
        RECT 5.330 882.585 494.230 885.415 ;
        RECT 5.330 877.145 494.230 879.975 ;
        RECT 5.330 871.705 494.230 874.535 ;
        RECT 5.330 866.265 494.230 869.095 ;
        RECT 5.330 860.825 494.230 863.655 ;
        RECT 5.330 855.385 494.230 858.215 ;
        RECT 5.330 849.945 494.230 852.775 ;
        RECT 5.330 844.505 494.230 847.335 ;
        RECT 5.330 839.065 494.230 841.895 ;
        RECT 5.330 833.625 494.230 836.455 ;
        RECT 5.330 828.185 494.230 831.015 ;
        RECT 5.330 822.745 494.230 825.575 ;
        RECT 5.330 817.305 494.230 820.135 ;
        RECT 5.330 811.865 494.230 814.695 ;
        RECT 5.330 806.425 494.230 809.255 ;
        RECT 5.330 800.985 494.230 803.815 ;
        RECT 5.330 795.545 494.230 798.375 ;
        RECT 5.330 790.105 494.230 792.935 ;
        RECT 5.330 784.665 494.230 787.495 ;
        RECT 5.330 779.225 494.230 782.055 ;
        RECT 5.330 773.785 494.230 776.615 ;
        RECT 5.330 768.345 494.230 771.175 ;
        RECT 5.330 762.905 494.230 765.735 ;
        RECT 5.330 757.465 494.230 760.295 ;
        RECT 5.330 752.025 494.230 754.855 ;
        RECT 5.330 746.585 494.230 749.415 ;
        RECT 5.330 741.145 494.230 743.975 ;
        RECT 5.330 735.705 494.230 738.535 ;
        RECT 5.330 730.265 494.230 733.095 ;
        RECT 5.330 724.825 494.230 727.655 ;
        RECT 5.330 719.385 494.230 722.215 ;
        RECT 5.330 713.945 494.230 716.775 ;
        RECT 5.330 708.505 494.230 711.335 ;
        RECT 5.330 703.065 494.230 705.895 ;
        RECT 5.330 697.625 494.230 700.455 ;
        RECT 5.330 692.185 494.230 695.015 ;
        RECT 5.330 686.745 494.230 689.575 ;
        RECT 5.330 681.305 494.230 684.135 ;
        RECT 5.330 675.865 494.230 678.695 ;
        RECT 5.330 670.425 494.230 673.255 ;
        RECT 5.330 664.985 494.230 667.815 ;
        RECT 5.330 659.545 494.230 662.375 ;
        RECT 5.330 654.105 494.230 656.935 ;
        RECT 5.330 648.665 494.230 651.495 ;
        RECT 5.330 643.225 494.230 646.055 ;
        RECT 5.330 637.785 494.230 640.615 ;
        RECT 5.330 632.345 494.230 635.175 ;
        RECT 5.330 626.905 494.230 629.735 ;
        RECT 5.330 621.465 494.230 624.295 ;
        RECT 5.330 616.025 494.230 618.855 ;
        RECT 5.330 610.585 494.230 613.415 ;
        RECT 5.330 605.145 494.230 607.975 ;
        RECT 5.330 599.705 494.230 602.535 ;
        RECT 5.330 594.265 494.230 597.095 ;
        RECT 5.330 588.825 494.230 591.655 ;
        RECT 5.330 583.385 494.230 586.215 ;
        RECT 5.330 577.945 494.230 580.775 ;
        RECT 5.330 572.505 494.230 575.335 ;
        RECT 5.330 567.065 494.230 569.895 ;
        RECT 5.330 561.625 494.230 564.455 ;
        RECT 5.330 556.185 494.230 559.015 ;
        RECT 5.330 550.745 494.230 553.575 ;
        RECT 5.330 545.305 494.230 548.135 ;
        RECT 5.330 539.865 494.230 542.695 ;
        RECT 5.330 534.425 494.230 537.255 ;
        RECT 5.330 528.985 494.230 531.815 ;
        RECT 5.330 523.545 494.230 526.375 ;
        RECT 5.330 518.105 494.230 520.935 ;
        RECT 5.330 512.665 494.230 515.495 ;
        RECT 5.330 507.225 494.230 510.055 ;
        RECT 5.330 501.785 494.230 504.615 ;
        RECT 5.330 496.345 494.230 499.175 ;
        RECT 5.330 490.905 494.230 493.735 ;
        RECT 5.330 485.465 494.230 488.295 ;
        RECT 5.330 480.025 494.230 482.855 ;
        RECT 5.330 474.585 494.230 477.415 ;
        RECT 5.330 469.145 494.230 471.975 ;
        RECT 5.330 463.705 494.230 466.535 ;
        RECT 5.330 458.265 494.230 461.095 ;
        RECT 5.330 452.825 494.230 455.655 ;
        RECT 5.330 447.385 494.230 450.215 ;
        RECT 5.330 441.945 494.230 444.775 ;
        RECT 5.330 436.505 494.230 439.335 ;
        RECT 5.330 431.065 494.230 433.895 ;
        RECT 5.330 425.625 494.230 428.455 ;
        RECT 5.330 420.185 494.230 423.015 ;
        RECT 5.330 414.745 494.230 417.575 ;
        RECT 5.330 409.305 494.230 412.135 ;
        RECT 5.330 403.865 494.230 406.695 ;
        RECT 5.330 398.425 494.230 401.255 ;
        RECT 5.330 392.985 494.230 395.815 ;
        RECT 5.330 387.545 494.230 390.375 ;
        RECT 5.330 382.105 494.230 384.935 ;
        RECT 5.330 376.665 494.230 379.495 ;
        RECT 5.330 371.225 494.230 374.055 ;
        RECT 5.330 365.785 494.230 368.615 ;
        RECT 5.330 360.345 494.230 363.175 ;
        RECT 5.330 354.905 494.230 357.735 ;
        RECT 5.330 349.465 494.230 352.295 ;
        RECT 5.330 344.025 494.230 346.855 ;
        RECT 5.330 338.585 494.230 341.415 ;
        RECT 5.330 333.145 494.230 335.975 ;
        RECT 5.330 327.705 494.230 330.535 ;
        RECT 5.330 322.265 494.230 325.095 ;
        RECT 5.330 316.825 494.230 319.655 ;
        RECT 5.330 311.385 494.230 314.215 ;
        RECT 5.330 305.945 494.230 308.775 ;
        RECT 5.330 300.505 494.230 303.335 ;
        RECT 5.330 295.065 494.230 297.895 ;
        RECT 5.330 289.625 494.230 292.455 ;
        RECT 5.330 284.185 494.230 287.015 ;
        RECT 5.330 278.745 494.230 281.575 ;
        RECT 5.330 273.305 494.230 276.135 ;
        RECT 5.330 267.865 494.230 270.695 ;
        RECT 5.330 262.425 494.230 265.255 ;
        RECT 5.330 256.985 494.230 259.815 ;
        RECT 5.330 251.545 494.230 254.375 ;
        RECT 5.330 246.105 494.230 248.935 ;
        RECT 5.330 240.665 494.230 243.495 ;
        RECT 5.330 235.225 494.230 238.055 ;
        RECT 5.330 229.785 494.230 232.615 ;
        RECT 5.330 224.345 494.230 227.175 ;
        RECT 5.330 218.905 494.230 221.735 ;
        RECT 5.330 213.465 494.230 216.295 ;
        RECT 5.330 208.025 494.230 210.855 ;
        RECT 5.330 202.585 494.230 205.415 ;
        RECT 5.330 197.145 494.230 199.975 ;
        RECT 5.330 191.705 494.230 194.535 ;
        RECT 5.330 186.265 494.230 189.095 ;
        RECT 5.330 180.825 494.230 183.655 ;
        RECT 5.330 175.385 494.230 178.215 ;
        RECT 5.330 169.945 494.230 172.775 ;
        RECT 5.330 164.505 494.230 167.335 ;
        RECT 5.330 159.065 494.230 161.895 ;
        RECT 5.330 153.625 494.230 156.455 ;
        RECT 5.330 148.185 494.230 151.015 ;
        RECT 5.330 142.745 494.230 145.575 ;
        RECT 5.330 137.305 494.230 140.135 ;
        RECT 5.330 131.865 494.230 134.695 ;
        RECT 5.330 126.425 494.230 129.255 ;
        RECT 5.330 120.985 494.230 123.815 ;
        RECT 5.330 115.545 494.230 118.375 ;
        RECT 5.330 110.105 494.230 112.935 ;
        RECT 5.330 104.665 494.230 107.495 ;
        RECT 5.330 99.225 494.230 102.055 ;
        RECT 5.330 93.785 494.230 96.615 ;
        RECT 5.330 88.345 494.230 91.175 ;
        RECT 5.330 82.905 494.230 85.735 ;
        RECT 5.330 77.465 494.230 80.295 ;
        RECT 5.330 72.025 494.230 74.855 ;
        RECT 5.330 66.585 494.230 69.415 ;
        RECT 5.330 61.145 494.230 63.975 ;
        RECT 5.330 55.705 494.230 58.535 ;
        RECT 5.330 50.265 494.230 53.095 ;
        RECT 5.330 44.825 494.230 47.655 ;
        RECT 5.330 39.385 494.230 42.215 ;
        RECT 5.330 33.945 494.230 36.775 ;
        RECT 5.330 28.505 494.230 31.335 ;
        RECT 5.330 23.065 494.230 25.895 ;
        RECT 5.330 17.625 494.230 20.455 ;
        RECT 5.330 12.185 494.230 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 494.040 2986.645 ;
      LAYER met1 ;
        RECT 5.520 10.640 494.040 2986.800 ;
      LAYER met2 ;
        RECT 12.150 2995.720 28.330 2996.490 ;
        RECT 29.170 2995.720 45.350 2996.490 ;
        RECT 46.190 2995.720 62.370 2996.490 ;
        RECT 63.210 2995.720 79.390 2996.490 ;
        RECT 80.230 2995.720 96.410 2996.490 ;
        RECT 97.250 2995.720 113.430 2996.490 ;
        RECT 114.270 2995.720 130.450 2996.490 ;
        RECT 131.290 2995.720 147.470 2996.490 ;
        RECT 148.310 2995.720 164.490 2996.490 ;
        RECT 165.330 2995.720 181.510 2996.490 ;
        RECT 182.350 2995.720 198.530 2996.490 ;
        RECT 199.370 2995.720 215.550 2996.490 ;
        RECT 216.390 2995.720 232.570 2996.490 ;
        RECT 233.410 2995.720 249.590 2996.490 ;
        RECT 250.430 2995.720 266.610 2996.490 ;
        RECT 267.450 2995.720 283.630 2996.490 ;
        RECT 284.470 2995.720 300.650 2996.490 ;
        RECT 301.490 2995.720 317.670 2996.490 ;
        RECT 318.510 2995.720 334.690 2996.490 ;
        RECT 335.530 2995.720 351.710 2996.490 ;
        RECT 352.550 2995.720 368.730 2996.490 ;
        RECT 369.570 2995.720 385.750 2996.490 ;
        RECT 386.590 2995.720 402.770 2996.490 ;
        RECT 403.610 2995.720 419.790 2996.490 ;
        RECT 420.630 2995.720 436.810 2996.490 ;
        RECT 437.650 2995.720 453.830 2996.490 ;
        RECT 454.670 2995.720 470.850 2996.490 ;
        RECT 471.690 2995.720 483.410 2996.490 ;
        RECT 11.870 4.280 483.410 2995.720 ;
        RECT 11.870 4.000 124.470 4.280 ;
        RECT 125.310 4.000 374.250 4.280 ;
        RECT 375.090 4.000 483.410 4.280 ;
      LAYER met3 ;
        RECT 21.050 10.715 483.430 2986.725 ;
  END
END user_proj_solar
END LIBRARY

